//----------------------------------------------------------------------------
// Task
//----------------------------------------------------------------------------

module formula_1_impl_2_fsm
(
    input               clk,
    input               rst,

    input               arg_vld,
    input        [31:0] a,
    input        [31:0] b,
    input        [31:0] c,

    output logic        res_vld,
    output logic [31:0] res,

    // isqrt interface

    output logic        isqrt_1_x_vld,
    output logic [31:0] isqrt_1_x,

    input               isqrt_1_y_vld,
    input        [15:0] isqrt_1_y,

    output logic        isqrt_2_x_vld,
    output logic [31:0] isqrt_2_x,

    input               isqrt_2_y_vld,
    input        [15:0] isqrt_2_y
);

    // Task:
    // Implement a module that calculates the folmula from the `formula_1_fn.svh` file
    // using two instances of the isqrt module in parallel.
    //
    // Design the FSM to calculate an answer and provide the correct `res` value    
    enum logic[1:0]
    {
      ST_IDLE        = 2'd0,
      ST_WAIT_RES_AB = 2'd1,
      ST_WAIT_RES_C  = 2'd2
    } state, next_state;

    always_comb begin
      next_state    = state;

      isqrt_1_x     = 'x;
      isqrt_1_x_vld = 1'b0;
      isqrt_2_x     = 'x;
      isqrt_2_x_vld = 1'b0;

      case(state)
        ST_IDLE: begin
	  isqrt_1_x = a;
	  isqrt_2_x = b;
	  if(arg_vld) begin
	    isqrt_1_x_vld = 1'b1;
	    isqrt_2_x_vld = 1'b1;
	    next_state    = ST_WAIT_RES_AB;
	  end
	end
	
        ST_WAIT_RES_AB: begin
	  isqrt_1_x = c;
	  isqrt_2_x = '0;
	  if(isqrt_1_y_vld && isqrt_2_y_vld) begin
	    isqrt_1_x_vld = 1'b1;
	    isqrt_2_x_vld = 1'b1;
	    next_state = ST_WAIT_RES_C;
	  end
	end

        ST_WAIT_RES_C: begin
	  if(isqrt_1_y_vld && isqrt_2_y_vld) begin
	    next_state = ST_IDLE;
	  end
	end
      endcase
    end

    always_ff @(posedge clk)
      if(rst)
        state <= ST_IDLE;
      else
	state <= next_state;

    always_ff @(posedge clk)
      if(state == ST_IDLE)
        res <= '0;
      else if(isqrt_1_y_vld && isqrt_2_y_vld)
	res <= res + isqrt_1_y + isqrt_2_y;

    always_ff @(posedge clk)
      if(rst)
	res_vld <= 1'b0;
      else
	res_vld <= (state == ST_WAIT_RES_C & (isqrt_1_y_vld & isqrt_2_y_vld));

endmodule
